module test (
  rstn,
  clk
);
input rstn;
input clk;

endmodule

